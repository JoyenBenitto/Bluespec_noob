// Making adder with funcitons instead of methods

package add;

    function int sum(int x, int y, int c);
    

endpackage: add