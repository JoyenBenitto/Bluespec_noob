package top

(*synthesize*)
module decode();


endmodule

endpackage